// Decode pipe bit positions
`define OPCODE_RANGE 6:0
`define FUNCT3_RANGE 9:7
`define FUNCT7_RANGE 16:10
`define RD_NUM_RANGE 21:17
`define OPERAND1_RANGE 53:22
`define OPERAND2_RANGE 85:54
`define OPERAND3_RANGE 117:86

`define DECODE_PIPE_MSB 117






// Execute pipe bit positions


`define EXECUTE_PIPE_MSB 8
