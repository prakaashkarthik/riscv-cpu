// Decode pipe bit positions
`define OPCODE_RANGE 6:0
`define FUNCT3_RANGE 9:7
`define RD_NUM_RANGE 14:10
`define RS1_NUM_RANGE 19:15
`define RS2_NUM_RANGE 24:20
`define RS1_DATA_RANGE 56:25
`define RS2_DATA_RANGE 88:57
`define IMM_DATA_RANGE 100:89

`define DECODE_PIPE_MSB 100
