localparam REGISTER_WIDTH = 32;

// Function specific register mnemnonics
`define ZERO 0
`define RA 1 // Return Address
`define SP 2 // Stack Pointer
`define GP 3 // Global Pointer
`define TP 4 // Thread Pointer
`define T0 5 // Temporary 0
`define T1 6 // Temporary 1
`define T2 7 // Temporary 2
`define FP 8 // Frame Pointer
`define S0 8 // Saved register 0
`define S1 9 // Saved register 1
`define A0 10 // Function argument / return value
`define A1 11 // Function argument / return value
`define A2 12 // Function argument
`define A3 13 
`define A4 14
`define A5 15
`define A6 16
`define A7 17
`define S2 18 // Saved register 2 - 11
`define S3 19
`define S4 20
`define S5 21
`define S6 22
`define S7 23
`define S8 24
`define S9 25
`define S10 26
`define S11 27
`define T3 28 // Temporary 3 - 6
`define T4 29
`define T5 30
`define T6 31

// Generic register mnemonics
`define X0 0
`define X1 1
`define X2 2
`define X3 3
`define X4 4
`define X5 5
`define X6 6
`define X7 7
`define X8 8
`define X9 9
`define X10 10
`define X11 11
`define X12 12
`define X13 13
`define X14 14
`define X15 15
`define X16 16
`define X17 17
`define X18 18
`define X19 19
`define X20 20
`define X21 21
`define X22 22
`define X23 23
`define X24 24
`define X25 25
`define X26 26
`define X27 27
`define X28 28
`define X29 29
`define X30 30
`define X31 31

